-- jtag_uart_sys_tb.vhd

-- Generated using ACDS version 13.0 156 at 2019.06.05.09:25:22

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jtag_uart_sys_tb is
end entity jtag_uart_sys_tb;

architecture rtl of jtag_uart_sys_tb is
	component jtag_uart_sys is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component jtag_uart_sys;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal jtag_uart_sys_inst_clk_bfm_clk_clk       : std_logic; -- jtag_uart_sys_inst_clk_bfm:clk -> [jtag_uart_sys_inst:clk_clk, jtag_uart_sys_inst_reset_bfm:clk]
	signal jtag_uart_sys_inst_reset_bfm_reset_reset : std_logic; -- jtag_uart_sys_inst_reset_bfm:reset -> jtag_uart_sys_inst:reset_reset_n

begin

	jtag_uart_sys_inst : component jtag_uart_sys
		port map (
			clk_clk       => jtag_uart_sys_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => jtag_uart_sys_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	jtag_uart_sys_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => jtag_uart_sys_inst_clk_bfm_clk_clk  -- clk.clk
		);

	jtag_uart_sys_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => jtag_uart_sys_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => jtag_uart_sys_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of jtag_uart_sys_tb
