library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity maquina_estados is
begin
end entity;

architecture arch of maquina_estados is

begin

end architecture;