// system_0.v

// Generated using ACDS version 13.0sp1 232 at 2019.07.17.12:55:16

`timescale 1 ps / 1 ps
module system_0 (
		input  wire        clk_50,                            //                   clk_50_clk_in.clk
		output wire [11:0] zs_addr_from_the_sdram_0,          //                    sdram_0_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram_0,            //                                .ba
		output wire        zs_cas_n_from_the_sdram_0,         //                                .cas_n
		output wire        zs_cke_from_the_sdram_0,           //                                .cke
		output wire        zs_cs_n_from_the_sdram_0,          //                                .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram_0,     //                                .dq
		output wire [1:0]  zs_dqm_from_the_sdram_0,           //                                .dqm
		output wire        zs_ras_n_from_the_sdram_0,         //                                .ras_n
		output wire        zs_we_n_from_the_sdram_0,          //                                .we_n
		inout  wire [7:0]  tri_state_bridge_0_data,           // tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		output wire [0:0]  tri_state_bridge_0_readn,          //                                .tri_state_bridge_0_readn
		output wire [0:0]  write_n_to_the_cfi_flash_0,        //                                .write_n_to_the_cfi_flash_0
		output wire [21:0] tri_state_bridge_0_address,        //                                .tri_state_bridge_0_address
		output wire [0:0]  select_n_to_the_cfi_flash_0,       //                                .select_n_to_the_cfi_flash_0
		input  wire        reset_n,                           //          merged_resets_in_reset.reset_n
		input  wire [3:0]  in_port_to_the_button_pio,         //  button_pio_external_connection.export
		input  wire [17:0] in_port_to_the_switch_pio,         //  switch_pio_external_connection.export
		input  wire        dm9000a_iOSC_50,                   //                         dm9000a.iOSC_50
		inout  wire [15:0] dm9000a_ENET_DATA,                 //                                .ENET_DATA
		output wire        dm9000a_ENET_CMD,                  //                                .ENET_CMD
		output wire        dm9000a_ENET_RD_N,                 //                                .ENET_RD_N
		output wire        dm9000a_ENET_WR_N,                 //                                .ENET_WR_N
		output wire        dm9000a_ENET_CS_N,                 //                                .ENET_CS_N
		output wire        dm9000a_ENET_RST_N,                //                                .ENET_RST_N
		output wire        dm9000a_ENET_CLK,                  //                                .ENET_CLK
		input  wire        dm9000a_ENET_INT,                  //                                .ENET_INT
		inout  wire [15:0] sram_0_avalon_slave_0_export_DQ,   //    sram_0_avalon_slave_0_export.DQ
		output wire [17:0] sram_0_avalon_slave_0_export_ADDR, //                                .ADDR
		output wire        sram_0_avalon_slave_0_export_UB_N, //                                .UB_N
		output wire        sram_0_avalon_slave_0_export_LB_N, //                                .LB_N
		output wire        sram_0_avalon_slave_0_export_WE_N, //                                .WE_N
		output wire        sram_0_avalon_slave_0_export_CE_N, //                                .CE_N
		output wire        sram_0_avalon_slave_0_export_OE_N, //                                .OE_N
		inout  wire        controller_pin_export              //                  controller_pin.export
	);

	wire    [0:0] tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out;                                        // tri_state_bridge_0_pinSharer_0:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_select_n_to_the_cfi_flash_0
	wire   [21:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out;                                         // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_address
	wire          tri_state_bridge_0_pinsharer_0_tcm_grant;                                                                  // tri_state_bridge_0_bridge_0:grant -> tri_state_bridge_0_pinSharer_0:grant
	wire    [0:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out;                                           // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_readn
	wire          tri_state_bridge_0_pinsharer_0_tcm_request;                                                                // tri_state_bridge_0_pinSharer_0:request -> tri_state_bridge_0_bridge_0:request
	wire    [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in;                                             // tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_in -> tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_in
	wire          tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen;                                          // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_outen -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_outen
	wire    [0:0] tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out;                                         // tri_state_bridge_0_pinSharer_0:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_write_n_to_the_cfi_flash_0
	wire    [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out;                                            // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data
	wire          cfi_flash_0_tcm_chipselect_n_out;                                                                          // cfi_flash_0:tcm_chipselect_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_chipselect_n_out
	wire          cfi_flash_0_tcm_grant;                                                                                     // tri_state_bridge_0_pinSharer_0:tcs0_grant -> cfi_flash_0:tcm_grant
	wire          cfi_flash_0_tcm_data_outen;                                                                                // cfi_flash_0:tcm_data_outen -> tri_state_bridge_0_pinSharer_0:tcs0_data_outen
	wire          cfi_flash_0_tcm_request;                                                                                   // cfi_flash_0:tcm_request -> tri_state_bridge_0_pinSharer_0:tcs0_request
	wire    [7:0] cfi_flash_0_tcm_data_out;                                                                                  // cfi_flash_0:tcm_data_out -> tri_state_bridge_0_pinSharer_0:tcs0_data_out
	wire          cfi_flash_0_tcm_write_n_out;                                                                               // cfi_flash_0:tcm_write_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_write_n_out
	wire   [21:0] cfi_flash_0_tcm_address_out;                                                                               // cfi_flash_0:tcm_address_out -> tri_state_bridge_0_pinSharer_0:tcs0_address_out
	wire    [7:0] cfi_flash_0_tcm_data_in;                                                                                   // tri_state_bridge_0_pinSharer_0:tcs0_data_in -> cfi_flash_0:tcm_data_in
	wire          cfi_flash_0_tcm_read_n_out;                                                                                // cfi_flash_0:tcm_read_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_read_n_out
	wire          cpu_0_instruction_master_waitrequest;                                                                      // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire   [24:0] cpu_0_instruction_master_address;                                                                          // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire          cpu_0_instruction_master_read;                                                                             // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire   [31:0] cpu_0_instruction_master_readdata;                                                                         // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire          cpu_0_data_master_waitrequest;                                                                             // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire   [31:0] cpu_0_data_master_writedata;                                                                               // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire   [24:0] cpu_0_data_master_address;                                                                                 // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire          cpu_0_data_master_write;                                                                                   // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire          cpu_0_data_master_read;                                                                                    // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire   [31:0] cpu_0_data_master_readdata;                                                                                // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire          cpu_0_data_master_debugaccess;                                                                             // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire    [3:0] cpu_0_data_master_byteenable;                                                                              // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                        // cpu_0:jtag_debug_module_waitrequest -> cpu_0_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                          // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire    [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                            // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                              // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                               // cpu_0_jtag_debug_module_translator:av_read -> cpu_0:jtag_debug_module_read
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                           // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire          cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                        // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire    [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                         // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire          sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                     // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                       // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire   [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                         // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire          sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                      // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire          sdram_0_s1_translator_avalon_anti_slave_0_write;                                                           // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire          sdram_0_s1_translator_avalon_anti_slave_0_read;                                                            // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                        // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire          sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                   // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire    [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                      // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire   [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata;                                // epcs_controller_epcs_control_port_translator:av_writedata -> epcs_controller:writedata
	wire    [8:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address;                                  // epcs_controller_epcs_control_port_translator:av_address -> epcs_controller:address
	wire          epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                               // epcs_controller_epcs_control_port_translator:av_chipselect -> epcs_controller:chipselect
	wire          epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write;                                    // epcs_controller_epcs_control_port_translator:av_write -> epcs_controller:write_n
	wire          epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read;                                     // epcs_controller_epcs_control_port_translator:av_read -> epcs_controller:read_n
	wire   [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata;                                 // epcs_controller:readdata -> epcs_controller_epcs_control_port_translator:av_readdata
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest;                                                // cfi_flash_0:uas_waitrequest -> cfi_flash_0_uas_translator:av_waitrequest
	wire    [0:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount;                                                 // cfi_flash_0_uas_translator:av_burstcount -> cfi_flash_0:uas_burstcount
	wire    [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata;                                                  // cfi_flash_0_uas_translator:av_writedata -> cfi_flash_0:uas_writedata
	wire   [21:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_address;                                                    // cfi_flash_0_uas_translator:av_address -> cfi_flash_0:uas_address
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_lock;                                                       // cfi_flash_0_uas_translator:av_lock -> cfi_flash_0:uas_lock
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_write;                                                      // cfi_flash_0_uas_translator:av_write -> cfi_flash_0:uas_write
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_read;                                                       // cfi_flash_0_uas_translator:av_read -> cfi_flash_0:uas_read
	wire    [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata;                                                   // cfi_flash_0:uas_readdata -> cfi_flash_0_uas_translator:av_readdata
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess;                                                // cfi_flash_0_uas_translator:av_debugaccess -> cfi_flash_0:uas_debugaccess
	wire          cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid;                                              // cfi_flash_0:uas_readdatavalid -> cfi_flash_0_uas_translator:av_readdatavalid
	wire    [0:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable;                                                 // cfi_flash_0_uas_translator:av_byteenable -> cfi_flash_0:uas_byteenable
	wire    [0:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                         // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                        // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                  // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                    // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                      // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                        // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                     // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                       // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire    [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                         // timer_0_s1_translator:av_address -> timer_0:address
	wire          timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                      // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire          timer_0_s1_translator_avalon_anti_slave_0_write;                                                           // timer_0_s1_translator:av_write -> timer_0:write_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                        // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                       // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire    [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                         // timer_1_s1_translator:av_address -> timer_1:address
	wire          timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                                      // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire          timer_1_s1_translator_avalon_anti_slave_0_write;                                                           // timer_1_s1_translator:av_write -> timer_1:write_n
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                        // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                    // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire    [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                      // button_pio_s1_translator:av_address -> button_pio:address
	wire          button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                   // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire          button_pio_s1_translator_avalon_anti_slave_0_write;                                                        // button_pio_s1_translator:av_write -> button_pio:write_n
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                     // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire    [1:0] switch_pio_s1_translator_avalon_anti_slave_0_address;                                                      // switch_pio_s1_translator:av_address -> switch_pio:address
	wire   [31:0] switch_pio_s1_translator_avalon_anti_slave_0_readdata;                                                     // switch_pio:readdata -> switch_pio_s1_translator:av_readdata
	wire   [15:0] dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                           // DM9000A_avalon_slave_0_translator:av_writedata -> DM9000A:iDATA
	wire    [0:0] dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address;                                             // DM9000A_avalon_slave_0_translator:av_address -> DM9000A:iCMD
	wire          dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                          // DM9000A_avalon_slave_0_translator:av_chipselect -> DM9000A:iCS_N
	wire          dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write;                                               // DM9000A_avalon_slave_0_translator:av_write -> DM9000A:iWR_N
	wire          dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                // DM9000A_avalon_slave_0_translator:av_read -> DM9000A:iRD_N
	wire   [15:0] dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                            // DM9000A:oDATA -> DM9000A_avalon_slave_0_translator:av_readdata
	wire   [15:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                            // sram_0_avalon_slave_0_translator:av_writedata -> sram_0:iDATA
	wire   [17:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                              // sram_0_avalon_slave_0_translator:av_address -> sram_0:iADDR
	wire          sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                           // sram_0_avalon_slave_0_translator:av_chipselect -> sram_0:iCE_N
	wire          sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                // sram_0_avalon_slave_0_translator:av_write -> sram_0:iWE_N
	wire          sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                                 // sram_0_avalon_slave_0_translator:av_read -> sram_0:iOE_N
	wire   [15:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                             // sram_0:oDATA -> sram_0_avalon_slave_0_translator:av_readdata
	wire    [1:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                           // sram_0_avalon_slave_0_translator:av_byteenable -> sram_0:iBE_N
	wire   [63:0] gamecube_controller_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // gamecube_controller_0:readdata -> gamecube_controller_0_avalon_slave_0_translator:av_readdata
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                                   // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                                     // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                        // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                       // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                        // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                                    // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                        // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                         // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                          // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [24:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                            // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_data_master_translator_avalon_universal_master_0_lock;                                               // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_data_master_translator_avalon_universal_master_0_write;                                              // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_data_master_translator_avalon_universal_master_0_read;                                               // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                           // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire          cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                        // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                         // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                      // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                            // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire   [24:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                             // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire   [24:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // epcs_controller_epcs_control_port_translator:uav_waitrequest -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_controller_epcs_control_port_translator:uav_burstcount
	wire   [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                  // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_controller_epcs_control_port_translator:uav_writedata
	wire   [24:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_controller_epcs_control_port_translator:uav_address
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                      // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_controller_epcs_control_port_translator:uav_write
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_controller_epcs_control_port_translator:uav_lock
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_controller_epcs_control_port_translator:uav_read
	wire   [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                   // epcs_controller_epcs_control_port_translator:uav_readdata -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // epcs_controller_epcs_control_port_translator:uav_readdatavalid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_controller_epcs_control_port_translator:uav_debugaccess
	wire    [3:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_controller_epcs_control_port_translator:uav_byteenable
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;               // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;               // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // cfi_flash_0_uas_translator:uav_waitrequest -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_0_uas_translator:uav_burstcount
	wire    [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_0_uas_translator:uav_writedata
	wire   [24:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_0_uas_translator:uav_address
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write;                                        // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_0_uas_translator:uav_write
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_0_uas_translator:uav_lock
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read;                                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_0_uas_translator:uav_read
	wire    [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // cfi_flash_0_uas_translator:uav_readdata -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // cfi_flash_0_uas_translator:uav_readdatavalid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_0_uas_translator:uav_debugaccess
	wire    [0:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_0_uas_translator:uav_byteenable
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [74:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [74:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire    [9:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire   [24:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [24:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire   [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire    [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire   [24:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire    [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire   [24:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire    [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // switch_pio_s1_translator:uav_waitrequest -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_pio_s1_translator:uav_burstcount
	wire   [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_pio_s1_translator:uav_writedata
	wire   [24:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_pio_s1_translator:uav_address
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_pio_s1_translator:uav_write
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_pio_s1_translator:uav_lock
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_pio_s1_translator:uav_read
	wire   [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // switch_pio_s1_translator:uav_readdata -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // switch_pio_s1_translator:uav_readdatavalid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_pio_s1_translator:uav_debugaccess
	wire    [3:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_pio_s1_translator:uav_byteenable
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // DM9000A_avalon_slave_0_translator:uav_waitrequest -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> DM9000A_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                             // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> DM9000A_avalon_slave_0_translator:uav_writedata
	wire   [24:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> DM9000A_avalon_slave_0_translator:uav_address
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                 // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> DM9000A_avalon_slave_0_translator:uav_write
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> DM9000A_avalon_slave_0_translator:uav_lock
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> DM9000A_avalon_slave_0_translator:uav_read
	wire   [31:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                              // DM9000A_avalon_slave_0_translator:uav_readdata -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // DM9000A_avalon_slave_0_translator:uav_readdatavalid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DM9000A_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> DM9000A_avalon_slave_0_translator:uav_byteenable
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                           // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // sram_0_avalon_slave_0_translator:uav_waitrequest -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_slave_0_translator:uav_burstcount
	wire   [15:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                              // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_slave_0_translator:uav_writedata
	wire   [24:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_slave_0_translator:uav_address
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                  // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_slave_0_translator:uav_write
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_slave_0_translator:uav_lock
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_slave_0_translator:uav_read
	wire   [15:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                               // sram_0_avalon_slave_0_translator:uav_readdata -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // sram_0_avalon_slave_0_translator:uav_readdatavalid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_slave_0_translator:uav_debugaccess
	wire    [1:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_slave_0_translator:uav_byteenable
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                            // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // gamecube_controller_0_avalon_slave_0_translator:uav_waitrequest -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [3:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> gamecube_controller_0_avalon_slave_0_translator:uav_burstcount
	wire   [63:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> gamecube_controller_0_avalon_slave_0_translator:uav_writedata
	wire   [24:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> gamecube_controller_0_avalon_slave_0_translator:uav_address
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> gamecube_controller_0_avalon_slave_0_translator:uav_write
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> gamecube_controller_0_avalon_slave_0_translator:uav_lock
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> gamecube_controller_0_avalon_slave_0_translator:uav_read
	wire   [63:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // gamecube_controller_0_avalon_slave_0_translator:uav_readdata -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // gamecube_controller_0_avalon_slave_0_translator:uav_readdatavalid -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gamecube_controller_0_avalon_slave_0_translator:uav_debugaccess
	wire    [7:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> gamecube_controller_0_avalon_slave_0_translator:uav_byteenable
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [137:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [137:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [65:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [100:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [100:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                      // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [100:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [82:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_001:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                      // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [100:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_002:sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                        // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [73:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data;                                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_003:sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [100:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_004:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [100:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_005:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [100:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_006:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [100:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_007:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [100:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_008:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [100:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_009:sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                 // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [100:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_010:sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                  // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [82:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_011:sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [136:0] gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_012:sink_ready -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                         // burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                               // burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                       // burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] burst_adapter_source0_data;                                                                                // burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [12:0] burst_adapter_source0_channel;                                                                             // burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                     // burst_adapter_001:source0_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                           // burst_adapter_001:source0_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                   // burst_adapter_001:source0_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [73:0] burst_adapter_001_source0_data;                                                                            // burst_adapter_001:source0_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [12:0] burst_adapter_001_source0_channel;                                                                         // burst_adapter_001:source0_channel -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                     // burst_adapter_002:source0_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                           // burst_adapter_002:source0_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                   // burst_adapter_002:source0_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] burst_adapter_002_source0_data;                                                                            // burst_adapter_002:source0_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                           // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [12:0] burst_adapter_002_source0_channel;                                                                         // burst_adapter_002:source0_channel -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cpu_0_jtag_debug_module_reset_reset;                                                                       // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                        // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cfi_flash_0:reset_reset, cfi_flash_0_uas_translator:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, epcs_controller:reset_n, epcs_controller_epcs_control_port_translator:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch_pio:reset_n, switch_pio_s1_translator:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tri_state_bridge_0_bridge_0:reset, tri_state_bridge_0_pinSharer_0:reset_reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_002_reset_out_reset;                                                                        // rst_controller_002:reset_out -> [DM9000A:iRST_N, DM9000A_avalon_slave_0_translator:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_002:reset, gamecube_controller_0:resetn, gamecube_controller_0_avalon_slave_0_translator:reset, gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, sram_0:iRST_N, sram_0_avalon_slave_0_translator:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                           // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                 // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                         // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src0_data;                                                                                  // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [12:0] cmd_xbar_demux_src0_channel;                                                                               // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                 // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                           // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                 // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                         // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src1_data;                                                                                  // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [12:0] cmd_xbar_demux_src1_channel;                                                                               // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                 // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                           // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                 // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                         // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src2_data;                                                                                  // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [12:0] cmd_xbar_demux_src2_channel;                                                                               // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                 // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                           // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                 // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                         // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src3_data;                                                                                  // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [12:0] cmd_xbar_demux_src3_channel;                                                                               // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                 // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                           // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                 // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                         // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src4_data;                                                                                  // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [12:0] cmd_xbar_demux_src4_channel;                                                                               // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                                 // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                       // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                             // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                     // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src0_data;                                                                              // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [12:0] cmd_xbar_demux_001_src0_channel;                                                                           // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                             // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                       // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                             // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                     // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src1_data;                                                                              // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [12:0] cmd_xbar_demux_001_src1_channel;                                                                           // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                             // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                       // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                             // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                     // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src2_data;                                                                              // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [12:0] cmd_xbar_demux_001_src2_channel;                                                                           // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                             // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                       // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                             // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                     // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src3_data;                                                                              // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [12:0] cmd_xbar_demux_001_src3_channel;                                                                           // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                             // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                       // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                             // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                     // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src4_data;                                                                              // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [12:0] cmd_xbar_demux_001_src4_channel;                                                                           // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                             // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                       // cmd_xbar_demux_001:src5_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                             // cmd_xbar_demux_001:src5_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                     // cmd_xbar_demux_001:src5_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src5_data;                                                                              // cmd_xbar_demux_001:src5_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src5_channel;                                                                           // cmd_xbar_demux_001:src5_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                       // cmd_xbar_demux_001:src6_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                             // cmd_xbar_demux_001:src6_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                     // cmd_xbar_demux_001:src6_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src6_data;                                                                              // cmd_xbar_demux_001:src6_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src6_channel;                                                                           // cmd_xbar_demux_001:src6_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                       // cmd_xbar_demux_001:src7_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                             // cmd_xbar_demux_001:src7_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                     // cmd_xbar_demux_001:src7_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src7_data;                                                                              // cmd_xbar_demux_001:src7_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src7_channel;                                                                           // cmd_xbar_demux_001:src7_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                       // cmd_xbar_demux_001:src8_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                             // cmd_xbar_demux_001:src8_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                     // cmd_xbar_demux_001:src8_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src8_data;                                                                              // cmd_xbar_demux_001:src8_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src8_channel;                                                                           // cmd_xbar_demux_001:src8_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                       // cmd_xbar_demux_001:src9_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                             // cmd_xbar_demux_001:src9_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                     // cmd_xbar_demux_001:src9_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src9_data;                                                                              // cmd_xbar_demux_001:src9_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src9_channel;                                                                           // cmd_xbar_demux_001:src9_channel -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                      // cmd_xbar_demux_001:src10_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                            // cmd_xbar_demux_001:src10_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                    // cmd_xbar_demux_001:src10_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src10_data;                                                                             // cmd_xbar_demux_001:src10_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_demux_001_src10_channel;                                                                          // cmd_xbar_demux_001:src10_channel -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                      // cmd_xbar_demux_001:src11_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                            // cmd_xbar_demux_001:src11_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                    // cmd_xbar_demux_001:src11_startofpacket -> width_adapter_004:in_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src11_data;                                                                             // cmd_xbar_demux_001:src11_data -> width_adapter_004:in_data
	wire   [12:0] cmd_xbar_demux_001_src11_channel;                                                                          // cmd_xbar_demux_001:src11_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                      // cmd_xbar_demux_001:src12_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                            // cmd_xbar_demux_001:src12_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                    // cmd_xbar_demux_001:src12_startofpacket -> width_adapter_006:in_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src12_data;                                                                             // cmd_xbar_demux_001:src12_data -> width_adapter_006:in_data
	wire   [12:0] cmd_xbar_demux_001_src12_channel;                                                                          // cmd_xbar_demux_001:src12_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                           // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                 // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                         // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src0_data;                                                                                  // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [12:0] rsp_xbar_demux_src0_channel;                                                                               // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                 // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                           // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                 // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                         // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src1_data;                                                                                  // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [12:0] rsp_xbar_demux_src1_channel;                                                                               // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                 // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                       // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                             // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                     // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src0_data;                                                                              // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [12:0] rsp_xbar_demux_001_src0_channel;                                                                           // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                             // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                       // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                             // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                     // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src1_data;                                                                              // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [12:0] rsp_xbar_demux_001_src1_channel;                                                                           // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                             // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                       // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                             // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                     // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [100:0] rsp_xbar_demux_002_src0_data;                                                                              // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [12:0] rsp_xbar_demux_002_src0_channel;                                                                           // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                             // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                       // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                             // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                     // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [100:0] rsp_xbar_demux_002_src1_data;                                                                              // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [12:0] rsp_xbar_demux_002_src1_channel;                                                                           // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                             // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                       // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                             // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                     // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [100:0] rsp_xbar_demux_003_src0_data;                                                                              // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [12:0] rsp_xbar_demux_003_src0_channel;                                                                           // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                             // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                       // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                             // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                     // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [100:0] rsp_xbar_demux_003_src1_data;                                                                              // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [12:0] rsp_xbar_demux_003_src1_channel;                                                                           // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                             // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                       // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                             // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                     // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [100:0] rsp_xbar_demux_004_src0_data;                                                                              // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [12:0] rsp_xbar_demux_004_src0_channel;                                                                           // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                             // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                       // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                             // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                     // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [100:0] rsp_xbar_demux_004_src1_data;                                                                              // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [12:0] rsp_xbar_demux_004_src1_channel;                                                                           // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                             // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                       // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                             // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                     // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [100:0] rsp_xbar_demux_005_src0_data;                                                                              // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [12:0] rsp_xbar_demux_005_src0_channel;                                                                           // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                             // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                       // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                             // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                     // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [100:0] rsp_xbar_demux_006_src0_data;                                                                              // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [12:0] rsp_xbar_demux_006_src0_channel;                                                                           // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                             // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                       // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                             // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                     // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [100:0] rsp_xbar_demux_007_src0_data;                                                                              // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [12:0] rsp_xbar_demux_007_src0_channel;                                                                           // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                             // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                       // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                             // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                     // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [100:0] rsp_xbar_demux_008_src0_data;                                                                              // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [12:0] rsp_xbar_demux_008_src0_channel;                                                                           // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                             // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                       // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                             // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                     // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [100:0] rsp_xbar_demux_009_src0_data;                                                                              // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [12:0] rsp_xbar_demux_009_src0_channel;                                                                           // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                             // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                       // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                             // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                     // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [100:0] rsp_xbar_demux_010_src0_data;                                                                              // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [12:0] rsp_xbar_demux_010_src0_channel;                                                                           // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                             // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                       // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                             // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                     // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [100:0] rsp_xbar_demux_011_src0_data;                                                                              // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [12:0] rsp_xbar_demux_011_src0_channel;                                                                           // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                             // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                       // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                             // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                     // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [100:0] rsp_xbar_demux_012_src0_data;                                                                              // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [12:0] rsp_xbar_demux_012_src0_channel;                                                                           // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                             // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          addr_router_src_endofpacket;                                                                               // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                     // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                             // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [100:0] addr_router_src_data;                                                                                      // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [12:0] addr_router_src_channel;                                                                                   // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                     // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                              // rsp_xbar_mux:src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                    // rsp_xbar_mux:src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                            // rsp_xbar_mux:src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_mux_src_data;                                                                                     // rsp_xbar_mux:src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [12:0] rsp_xbar_mux_src_channel;                                                                                  // rsp_xbar_mux:src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                    // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                           // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                 // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                         // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [100:0] addr_router_001_src_data;                                                                                  // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [12:0] addr_router_001_src_channel;                                                                               // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                 // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                          // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                        // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_mux_001_src_data;                                                                                 // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [12:0] rsp_xbar_mux_001_src_channel;                                                                              // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                              // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                    // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                            // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_src_data;                                                                                     // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_mux_src_channel;                                                                                  // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                 // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                       // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                               // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [100:0] id_router_src_data;                                                                                        // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [12:0] id_router_src_channel;                                                                                     // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                       // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                          // cmd_xbar_mux_002:src_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                // cmd_xbar_mux_002:src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                        // cmd_xbar_mux_002:src_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_002_src_data;                                                                                 // cmd_xbar_mux_002:src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_mux_002_src_channel;                                                                              // cmd_xbar_mux_002:src_channel -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                             // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                   // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                           // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [100:0] id_router_002_src_data;                                                                                    // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [12:0] id_router_002_src_channel;                                                                                 // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                   // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                          // cmd_xbar_mux_004:src_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                                // cmd_xbar_mux_004:src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                        // cmd_xbar_mux_004:src_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_004_src_data;                                                                                 // cmd_xbar_mux_004:src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [12:0] cmd_xbar_mux_004_src_channel;                                                                              // cmd_xbar_mux_004:src_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                             // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                   // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                           // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [100:0] id_router_004_src_data;                                                                                    // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [12:0] id_router_004_src_channel;                                                                                 // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                   // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                             // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                   // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                           // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [100:0] id_router_005_src_data;                                                                                    // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [12:0] id_router_005_src_channel;                                                                                 // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                   // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                             // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                             // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                   // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                           // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [100:0] id_router_006_src_data;                                                                                    // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [12:0] id_router_006_src_channel;                                                                                 // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                   // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                             // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                             // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                   // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                           // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [100:0] id_router_007_src_data;                                                                                    // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [12:0] id_router_007_src_channel;                                                                                 // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                   // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                             // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                             // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                   // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                           // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [100:0] id_router_008_src_data;                                                                                    // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [12:0] id_router_008_src_channel;                                                                                 // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                   // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                             // switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                             // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                   // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                           // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [100:0] id_router_009_src_data;                                                                                    // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [12:0] id_router_009_src_channel;                                                                                 // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                   // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                            // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                             // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                   // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                           // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [100:0] id_router_010_src_data;                                                                                    // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [12:0] id_router_010_src_channel;                                                                                 // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                   // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                          // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                        // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [100:0] cmd_xbar_mux_001_src_data;                                                                                 // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [12:0] cmd_xbar_mux_001_src_channel;                                                                              // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                             // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                   // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                           // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [82:0] width_adapter_src_data;                                                                                    // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                   // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [12:0] width_adapter_src_channel;                                                                                 // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                             // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                                   // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                           // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [82:0] id_router_001_src_data;                                                                                    // id_router_001:src_data -> width_adapter_001:in_data
	wire   [12:0] id_router_001_src_channel;                                                                                 // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                                   // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                         // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                               // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                       // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [100:0] width_adapter_001_src_data;                                                                                // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                               // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [12:0] width_adapter_001_src_channel;                                                                             // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                          // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                        // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [100:0] cmd_xbar_mux_003_src_data;                                                                                 // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire   [12:0] cmd_xbar_mux_003_src_channel;                                                                              // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                         // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                               // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                       // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [73:0] width_adapter_002_src_data;                                                                                // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                               // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [12:0] width_adapter_002_src_channel;                                                                             // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_003_src_endofpacket;                                                                             // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_003_src_valid;                                                                                   // id_router_003:src_valid -> width_adapter_003:in_valid
	wire          id_router_003_src_startofpacket;                                                                           // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [73:0] id_router_003_src_data;                                                                                    // id_router_003:src_data -> width_adapter_003:in_data
	wire   [12:0] id_router_003_src_channel;                                                                                 // id_router_003:src_channel -> width_adapter_003:in_channel
	wire          id_router_003_src_ready;                                                                                   // width_adapter_003:in_ready -> id_router_003:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                         // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                               // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                       // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [100:0] width_adapter_003_src_data;                                                                                // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire          width_adapter_003_src_ready;                                                                               // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire   [12:0] width_adapter_003_src_channel;                                                                             // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                            // width_adapter_004:in_ready -> cmd_xbar_demux_001:src11_ready
	wire          width_adapter_004_src_endofpacket;                                                                         // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                               // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                       // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [82:0] width_adapter_004_src_data;                                                                                // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire          width_adapter_004_src_ready;                                                                               // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire   [12:0] width_adapter_004_src_channel;                                                                             // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire          id_router_011_src_endofpacket;                                                                             // id_router_011:src_endofpacket -> width_adapter_005:in_endofpacket
	wire          id_router_011_src_valid;                                                                                   // id_router_011:src_valid -> width_adapter_005:in_valid
	wire          id_router_011_src_startofpacket;                                                                           // id_router_011:src_startofpacket -> width_adapter_005:in_startofpacket
	wire   [82:0] id_router_011_src_data;                                                                                    // id_router_011:src_data -> width_adapter_005:in_data
	wire   [12:0] id_router_011_src_channel;                                                                                 // id_router_011:src_channel -> width_adapter_005:in_channel
	wire          id_router_011_src_ready;                                                                                   // width_adapter_005:in_ready -> id_router_011:src_ready
	wire          width_adapter_005_src_endofpacket;                                                                         // width_adapter_005:out_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          width_adapter_005_src_valid;                                                                               // width_adapter_005:out_valid -> rsp_xbar_demux_011:sink_valid
	wire          width_adapter_005_src_startofpacket;                                                                       // width_adapter_005:out_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [100:0] width_adapter_005_src_data;                                                                                // width_adapter_005:out_data -> rsp_xbar_demux_011:sink_data
	wire          width_adapter_005_src_ready;                                                                               // rsp_xbar_demux_011:sink_ready -> width_adapter_005:out_ready
	wire   [12:0] width_adapter_005_src_channel;                                                                             // width_adapter_005:out_channel -> rsp_xbar_demux_011:sink_channel
	wire          cmd_xbar_demux_001_src12_ready;                                                                            // width_adapter_006:in_ready -> cmd_xbar_demux_001:src12_ready
	wire          width_adapter_006_src_endofpacket;                                                                         // width_adapter_006:out_endofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_006_src_valid;                                                                               // width_adapter_006:out_valid -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_006_src_startofpacket;                                                                       // width_adapter_006:out_startofpacket -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [136:0] width_adapter_006_src_data;                                                                                // width_adapter_006:out_data -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_006_src_ready;                                                                               // gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_006:out_ready
	wire   [12:0] width_adapter_006_src_channel;                                                                             // width_adapter_006:out_channel -> gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_012_src_endofpacket;                                                                             // id_router_012:src_endofpacket -> width_adapter_007:in_endofpacket
	wire          id_router_012_src_valid;                                                                                   // id_router_012:src_valid -> width_adapter_007:in_valid
	wire          id_router_012_src_startofpacket;                                                                           // id_router_012:src_startofpacket -> width_adapter_007:in_startofpacket
	wire  [136:0] id_router_012_src_data;                                                                                    // id_router_012:src_data -> width_adapter_007:in_data
	wire   [12:0] id_router_012_src_channel;                                                                                 // id_router_012:src_channel -> width_adapter_007:in_channel
	wire          id_router_012_src_ready;                                                                                   // width_adapter_007:in_ready -> id_router_012:src_ready
	wire          width_adapter_007_src_endofpacket;                                                                         // width_adapter_007:out_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          width_adapter_007_src_valid;                                                                               // width_adapter_007:out_valid -> rsp_xbar_demux_012:sink_valid
	wire          width_adapter_007_src_startofpacket;                                                                       // width_adapter_007:out_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [100:0] width_adapter_007_src_data;                                                                                // width_adapter_007:out_data -> rsp_xbar_demux_012:sink_data
	wire          width_adapter_007_src_ready;                                                                               // rsp_xbar_demux_012:sink_ready -> width_adapter_007:out_ready
	wire   [12:0] width_adapter_007_src_channel;                                                                             // width_adapter_007:out_channel -> rsp_xbar_demux_012:sink_channel
	wire          irq_mapper_receiver0_irq;                                                                                  // epcs_controller:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                  // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                  // timer_0:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                  // timer_1:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                  // button_pio:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                  // DM9000A:oINT -> irq_mapper:receiver5_irq
	wire   [31:0] cpu_0_d_irq_irq;                                                                                           // irq_mapper:sender_irq -> cpu_0:d_irq

	system_0_sdram_0 sdram_0 (
		.clk            (clk_50),                                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                     // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram_0),                                //  wire.export
		.zs_ba          (zs_ba_from_the_sdram_0),                                  //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram_0),                               //      .export
		.zs_cke         (zs_cke_from_the_sdram_0),                                 //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram_0),                                //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram_0),                           //      .export
		.zs_dqm         (zs_dqm_from_the_sdram_0),                                 //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram_0),                               //      .export
		.zs_we_n        (zs_we_n_from_the_sdram_0)                                 //      .export
	);

	system_0_epcs_controller epcs_controller (
		.clk           (clk_50),                                                                      //               clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                         //             reset.reset_n
		.address       (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                            //                  .dataavailable
		.endofpacket   (),                                                                            //                  .endofpacket
		.read_n        (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                            //                  .readyfordata
		.write_n       (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq)                                                     //               irq.irq
	);

	system_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_50),                                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	system_0_timer_0 timer_0 (
		.clk        (clk_50),                                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                              //   irq.irq
	);

	system_0_timer_0 timer_1 (
		.clk        (clk_50),                                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                              //   irq.irq
	);

	system_0_button_pio button_pio (
		.clk        (clk_50),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_button_pio),                               // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                                 //                 irq.irq
	);

	system_0_switch_pio switch_pio (
		.clk      (clk_50),                                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address  (switch_pio_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_pio_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_switch_pio)                              // external_connection.export
	);

	system_0_cpu_0 cpu_0 (
		.clk                                   (clk_50),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	system_0_tri_state_bridge_0_bridge_0 tri_state_bridge_0_bridge_0 (
		.clk                               (clk_50),                                                             //   clk.clk
		.reset                             (rst_controller_001_reset_out_reset),                                 // reset.reset
		.request                           (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcs.request
		.grant                             (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tcs_tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tcs_tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.tcs_tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tcs_tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.tcs_write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tcs_tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tcs_select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data           (tri_state_bridge_0_data),                                            //   out.tri_state_bridge_0_data
		.tri_state_bridge_0_readn          (tri_state_bridge_0_readn),                                           //      .tri_state_bridge_0_readn
		.write_n_to_the_cfi_flash_0        (write_n_to_the_cfi_flash_0),                                         //      .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_address        (tri_state_bridge_0_address),                                         //      .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0       (select_n_to_the_cfi_flash_0)                                         //      .select_n_to_the_cfi_flash_0
	);

	system_0_tri_state_bridge_0_pinSharer_0 tri_state_bridge_0_pinsharer_0 (
		.clk_clk                       (clk_50),                                                             //   clk.clk
		.reset_reset                   (rst_controller_001_reset_out_reset),                                 // reset.reset
		.request                       (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcm.request
		.grant                         (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tcs0_request                  (cfi_flash_0_tcm_request),                                            //  tcs0.request
		.tcs0_grant                    (cfi_flash_0_tcm_grant),                                              //      .grant
		.tcs0_address_out              (cfi_flash_0_tcm_address_out),                                        //      .address_out
		.tcs0_read_n_out               (cfi_flash_0_tcm_read_n_out),                                         //      .read_n_out
		.tcs0_write_n_out              (cfi_flash_0_tcm_write_n_out),                                        //      .write_n_out
		.tcs0_data_out                 (cfi_flash_0_tcm_data_out),                                           //      .data_out
		.tcs0_data_in                  (cfi_flash_0_tcm_data_in),                                            //      .data_in
		.tcs0_data_outen               (cfi_flash_0_tcm_data_outen),                                         //      .data_outen
		.tcs0_chipselect_n_out         (cfi_flash_0_tcm_chipselect_n_out)                                    //      .chipselect_n_out
	);

	system_0_cfi_flash_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash_0 (
		.clk_clk              (clk_50),                                                       //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                           // reset.reset
		.uas_address          (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_0_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_0_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_0_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (cfi_flash_0_tcm_request),                                      //      .request
		.tcm_grant            (cfi_flash_0_tcm_grant),                                        //      .grant
		.tcm_address_out      (cfi_flash_0_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (cfi_flash_0_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (cfi_flash_0_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (cfi_flash_0_tcm_data_in)                                       //      .data_in
	);

	system_0_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_50),                                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                                //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	DM9000A_IF dm9000a (
		.iCLK       (clk_50),                                                            //                   clk.clk
		.iRST_N     (~rst_controller_002_reset_out_reset),                               //             clk_reset.reset_n
		.iOSC_50    (dm9000a_iOSC_50),                                                   // avalon_slave_0_export.export
		.ENET_DATA  (dm9000a_ENET_DATA),                                                 //                      .export
		.ENET_CMD   (dm9000a_ENET_CMD),                                                  //                      .export
		.ENET_RD_N  (dm9000a_ENET_RD_N),                                                 //                      .export
		.ENET_WR_N  (dm9000a_ENET_WR_N),                                                 //                      .export
		.ENET_CS_N  (dm9000a_ENET_CS_N),                                                 //                      .export
		.ENET_RST_N (dm9000a_ENET_RST_N),                                                //                      .export
		.ENET_CLK   (dm9000a_ENET_CLK),                                                  //                      .export
		.ENET_INT   (dm9000a_ENET_INT),                                                  //                      .export
		.iDATA      (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //        avalon_slave_0.writedata
		.iCMD       (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                      .address
		.iRD_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read_n
		.iWR_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write_n
		.iCS_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect_n
		.oDATA      (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                      .readdata
		.oINT       (irq_mapper_receiver5_irq)                                           //    avalon_slave_0_irq.irq
	);

	SRAM_16Bit_512K sram_0 (
		.iCLK      (clk_50),                                                           //                   clk.clk
		.iRST_N    (~rst_controller_002_reset_out_reset),                              //             clk_reset.reset_n
		.SRAM_DQ   (sram_0_avalon_slave_0_export_DQ),                                  // avalon_slave_0_export.export
		.SRAM_ADDR (sram_0_avalon_slave_0_export_ADDR),                                //                      .export
		.SRAM_UB_N (sram_0_avalon_slave_0_export_UB_N),                                //                      .export
		.SRAM_LB_N (sram_0_avalon_slave_0_export_LB_N),                                //                      .export
		.SRAM_WE_N (sram_0_avalon_slave_0_export_WE_N),                                //                      .export
		.SRAM_CE_N (sram_0_avalon_slave_0_export_CE_N),                                //                      .export
		.SRAM_OE_N (sram_0_avalon_slave_0_export_OE_N),                                //                      .export
		.iDATA     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //        avalon_slave_0.writedata
		.oDATA     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                      .readdata
		.iADDR     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                      .address
		.iWE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write_n
		.iOE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read_n
		.iCE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect_n
		.iBE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable)  //                      .byteenable_n
	);

	gc_avalon_interface gamecube_controller_0 (
		.readdata (gamecube_controller_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata), // avalon_slave_0.readdata
		.ctrl_pin (controller_pin_export),                                                        //    conduit_end.export
		.clock    (clk_50),                                                                       //     clock_sink.clk
		.resetn   (~rst_controller_002_reset_out_reset)                                           //     reset_sink.reset_n
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                      (clk_50),                                                                      //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address              (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_0_data_master_translator (
		.clk                      (clk_50),                                                               //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                     reset.reset
		.uav_address              (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_0_data_master_read),                                               //                          .read
		.av_readdata              (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_0_data_master_write),                                              //                          .write
		.av_writedata             (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                      (clk_50),                                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                      (clk_50),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_controller_epcs_control_port_translator (
		.clk                      (clk_50),                                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                             //              (terminated)
		.av_byteenable            (),                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                             //              (terminated)
		.av_lock                  (),                                                                                             //              (terminated)
		.av_clken                 (),                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                             //              (terminated)
		.uav_response             (),                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cfi_flash_0_uas_translator (
		.clk                      (clk_50),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock                  (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess           (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                      (clk_50),                                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                                      //              (terminated)
		.av_read                  (),                                                                                      //              (terminated)
		.av_writedata             (),                                                                                      //              (terminated)
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_byteenable            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_50),                                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (clk_50),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                      (clk_50),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                      (clk_50),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_pio_s1_translator (
		.clk                      (clk_50),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (switch_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                         //              (terminated)
		.av_read                  (),                                                                         //              (terminated)
		.av_writedata             (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dm9000a_avalon_slave_0_translator (
		.clk                      (clk_50),                                                                            //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                //                    reset.reset
		.uav_address              (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (1)
	) sram_0_avalon_slave_0_translator (
		.clk                      (clk_50),                                                                           //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                               //                    reset.reset
		.uav_address              (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) gamecube_controller_0_avalon_slave_0_translator (
		.clk                      (clk_50),                                                                                          //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                              //                    reset.reset
		.uav_address              (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_readdata              (gamecube_controller_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //      avalon_anti_slave_0.readdata
		.av_address               (),                                                                                                //              (terminated)
		.av_write                 (),                                                                                                //              (terminated)
		.av_read                  (),                                                                                                //              (terminated)
		.av_writedata             (),                                                                                                //              (terminated)
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_byteenable            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_chipselect            (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_50),                                                                               //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                               //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_50),                                                                        //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.av_address              (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                   //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                           //                .channel
		.rf_sink_ready           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (56),
		.PKT_DEST_ID_H             (63),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (46),
		.PKT_BURSTWRAP_L           (44),
		.PKT_BYTE_CNT_H            (43),
		.PKT_BYTE_CNT_L            (40),
		.PKT_PROTECTION_H          (67),
		.PKT_PROTECTION_L          (65),
		.PKT_RESPONSE_STATUS_H     (73),
		.PKT_RESPONSE_STATUS_L     (72),
		.PKT_BURST_SIZE_H          (49),
		.PKT_BURST_SIZE_L          (47),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (74),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                      //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                      //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                       //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                    //                .channel
		.rf_sink_ready           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (75),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (10),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_50),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                           // (terminated)
		.out_startofpacket (),                                                                               // (terminated)
		.out_endofpacket   (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                                    //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                 //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                    //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                    //                .channel
		.rf_sink_ready           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                      //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                            //                .channel
		.rf_sink_ready           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                     //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                          //                .channel
		.rf_sink_ready           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                     //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (117),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (96),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (97),
		.PKT_TRANS_POSTED          (98),
		.PKT_TRANS_WRITE           (99),
		.PKT_TRANS_READ            (100),
		.PKT_TRANS_LOCK            (101),
		.PKT_SRC_ID_H              (122),
		.PKT_SRC_ID_L              (119),
		.PKT_DEST_ID_H             (126),
		.PKT_DEST_ID_L             (123),
		.PKT_BURSTWRAP_H           (109),
		.PKT_BURSTWRAP_L           (107),
		.PKT_BYTE_CNT_H            (106),
		.PKT_BYTE_CNT_L            (103),
		.PKT_PROTECTION_H          (130),
		.PKT_PROTECTION_L          (128),
		.PKT_RESPONSE_STATUS_H     (136),
		.PKT_RESPONSE_STATUS_L     (135),
		.PKT_BURST_SIZE_H          (112),
		.PKT_BURST_SIZE_L          (110),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (137),
		.AVS_BURSTCOUNT_W          (4),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50),                                                                                                    //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_006_src_ready),                                                                               //              cp.ready
		.cp_valid                (width_adapter_006_src_valid),                                                                               //                .valid
		.cp_data                 (width_adapter_006_src_data),                                                                                //                .data
		.cp_startofpacket        (width_adapter_006_src_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (width_adapter_006_src_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (width_adapter_006_src_channel),                                                                             //                .channel
		.rf_sink_ready           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (138),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50),                                                                                                    //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	system_0_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	system_0_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	system_0_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	system_0_id_router_001 id_router_001 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                               //       src.ready
		.src_valid          (id_router_001_src_valid),                                               //          .valid
		.src_data           (id_router_001_src_data),                                                //          .data
		.src_channel        (id_router_001_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router id_router_002 (
		.sink_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                      //          .valid
		.src_data           (id_router_002_src_data),                                                                       //          .data
		.src_channel        (id_router_002_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                                 //          .endofpacket
	);

	system_0_id_router_003 id_router_003 (
		.sink_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                    //       src.ready
		.src_valid          (id_router_003_src_valid),                                                    //          .valid
		.src_data           (id_router_003_src_data),                                                     //          .data
		.src_channel        (id_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                               //          .endofpacket
	);

	system_0_id_router id_router_004 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                                               //          .valid
		.src_data           (id_router_004_src_data),                                                                //          .data
		.src_channel        (id_router_004_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_005 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	system_0_id_router_005 id_router_006 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_007 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                               //          .valid
		.src_data           (id_router_007_src_data),                                                //          .data
		.src_channel        (id_router_007_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_008 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                  //       src.ready
		.src_valid          (id_router_008_src_valid),                                                  //          .valid
		.src_data           (id_router_008_src_data),                                                   //          .data
		.src_channel        (id_router_008_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_005 id_router_009 (
		.sink_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                  //       src.ready
		.src_valid          (id_router_009_src_valid),                                                  //          .valid
		.src_data           (id_router_009_src_data),                                                   //          .data
		.src_channel        (id_router_009_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_005 id_router_010 (
		.sink_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                           //       src.ready
		.src_valid          (id_router_010_src_valid),                                                           //          .valid
		.src_data           (id_router_010_src_data),                                                            //          .data
		.src_channel        (id_router_010_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                      //          .endofpacket
	);

	system_0_id_router_011 id_router_011 (
		.sink_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                          //       src.ready
		.src_valid          (id_router_011_src_valid),                                                          //          .valid
		.src_data           (id_router_011_src_data),                                                           //          .data
		.src_channel        (id_router_011_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                     //          .endofpacket
	);

	system_0_id_router_012 id_router_012 (
		.sink_ready         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (gamecube_controller_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50),                                                                                          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_012_src_valid),                                                                         //          .valid
		.src_data           (id_router_012_src_data),                                                                          //          .data
		.src_channel        (id_router_012_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                                    //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (63),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (13),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (55),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_50),                              //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (43),
		.PKT_BYTE_CNT_L            (40),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (49),
		.PKT_BURST_SIZE_L          (47),
		.PKT_BURST_TYPE_H          (51),
		.PKT_BURST_TYPE_L          (50),
		.PKT_BURSTWRAP_H           (46),
		.PKT_BURSTWRAP_L           (44),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (74),
		.ST_CHANNEL_W              (13),
		.OUT_BYTE_CNT_H            (40),
		.OUT_BURSTWRAP_H           (46),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (clk_50),                                  //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (63),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (13),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (55),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clk_50),                                  //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (),                                    //       clk.clk
		.reset_out  (),                                    // reset_out.reset
		.reset_req  (),                                    // (terminated)
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (cpu_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.clk        (clk_50),                              //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req  (),                                    // (terminated)
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (clk_50),                             //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	system_0_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_50),                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),    //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),          //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),          //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),           //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),        //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)     //          .endofpacket
	);

	system_0_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_50),                                 //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_50),                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_007 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_008 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_009 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_012 (
		.clk                (clk_50),                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_007_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_007_src_channel),         //          .channel
		.sink_data          (width_adapter_007_src_data),            //          .data
		.sink_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_007_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_50),                                //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_50),                                //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (100),
		.IN_PKT_RESPONSE_STATUS_L      (99),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (101),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (52),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (58),
		.OUT_PKT_BURST_SIZE_L          (56),
		.OUT_PKT_RESPONSE_STATUS_H     (82),
		.OUT_PKT_RESPONSE_STATUS_L     (81),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (60),
		.OUT_PKT_BURST_TYPE_L          (59),
		.OUT_ST_DATA_W                 (83),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_50),                             //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (52),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (55),
		.IN_PKT_BURSTWRAP_L            (53),
		.IN_PKT_BURST_SIZE_H           (58),
		.IN_PKT_BURST_SIZE_L           (56),
		.IN_PKT_RESPONSE_STATUS_H      (82),
		.IN_PKT_RESPONSE_STATUS_L      (81),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (60),
		.IN_PKT_BURST_TYPE_L           (59),
		.IN_ST_DATA_W                  (83),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (100),
		.OUT_PKT_RESPONSE_STATUS_L     (99),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (101),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (100),
		.IN_PKT_RESPONSE_STATUS_L      (99),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (101),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (43),
		.OUT_PKT_BYTE_CNT_L            (40),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_PKT_BURST_SIZE_H          (49),
		.OUT_PKT_BURST_SIZE_L          (47),
		.OUT_PKT_RESPONSE_STATUS_H     (73),
		.OUT_PKT_RESPONSE_STATUS_L     (72),
		.OUT_PKT_TRANS_EXCLUSIVE       (39),
		.OUT_PKT_BURST_TYPE_H          (51),
		.OUT_PKT_BURST_TYPE_L          (50),
		.OUT_ST_DATA_W                 (74),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (43),
		.IN_PKT_BYTE_CNT_L             (40),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (46),
		.IN_PKT_BURSTWRAP_L            (44),
		.IN_PKT_BURST_SIZE_H           (49),
		.IN_PKT_BURST_SIZE_L           (47),
		.IN_PKT_RESPONSE_STATUS_H      (73),
		.IN_PKT_RESPONSE_STATUS_L      (72),
		.IN_PKT_TRANS_EXCLUSIVE        (39),
		.IN_PKT_BURST_TYPE_H           (51),
		.IN_PKT_BURST_TYPE_L           (50),
		.IN_ST_DATA_W                  (74),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (100),
		.OUT_PKT_RESPONSE_STATUS_L     (99),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (101),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_003_src_valid),             //      sink.valid
		.in_channel           (id_router_003_src_channel),           //          .channel
		.in_startofpacket     (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_003_src_ready),             //          .ready
		.in_data              (id_router_003_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (100),
		.IN_PKT_RESPONSE_STATUS_L      (99),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (101),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (52),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (58),
		.OUT_PKT_BURST_SIZE_L          (56),
		.OUT_PKT_RESPONSE_STATUS_H     (82),
		.OUT_PKT_RESPONSE_STATUS_L     (81),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (60),
		.OUT_PKT_BURST_TYPE_L          (59),
		.OUT_ST_DATA_W                 (83),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (clk_50),                                 //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src11_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src11_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src11_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src11_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (52),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (55),
		.IN_PKT_BURSTWRAP_L            (53),
		.IN_PKT_BURST_SIZE_H           (58),
		.IN_PKT_BURST_SIZE_L           (56),
		.IN_PKT_RESPONSE_STATUS_H      (82),
		.IN_PKT_RESPONSE_STATUS_L      (81),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (60),
		.IN_PKT_BURST_TYPE_L           (59),
		.IN_ST_DATA_W                  (83),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (100),
		.OUT_PKT_RESPONSE_STATUS_L     (99),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (101),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_011_src_valid),             //      sink.valid
		.in_channel           (id_router_011_src_channel),           //          .channel
		.in_startofpacket     (id_router_011_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_011_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_011_src_ready),             //          .ready
		.in_data              (id_router_011_src_data),              //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_005_src_data),          //          .data
		.out_channel          (width_adapter_005_src_channel),       //          .channel
		.out_valid            (width_adapter_005_src_valid),         //          .valid
		.out_ready            (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (100),
		.IN_PKT_RESPONSE_STATUS_L      (99),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (101),
		.OUT_PKT_ADDR_H                (96),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (106),
		.OUT_PKT_BYTE_CNT_L            (103),
		.OUT_PKT_TRANS_COMPRESSED_READ (97),
		.OUT_PKT_BURST_SIZE_H          (112),
		.OUT_PKT_BURST_SIZE_L          (110),
		.OUT_PKT_RESPONSE_STATUS_H     (136),
		.OUT_PKT_RESPONSE_STATUS_L     (135),
		.OUT_PKT_TRANS_EXCLUSIVE       (102),
		.OUT_PKT_BURST_TYPE_H          (114),
		.OUT_PKT_BURST_TYPE_L          (113),
		.OUT_ST_DATA_W                 (137),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_006 (
		.clk                  (clk_50),                                 //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src12_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src12_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src12_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src12_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_006_src_data),             //          .data
		.out_channel          (width_adapter_006_src_channel),          //          .channel
		.out_valid            (width_adapter_006_src_valid),            //          .valid
		.out_ready            (width_adapter_006_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (96),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (106),
		.IN_PKT_BYTE_CNT_L             (103),
		.IN_PKT_TRANS_COMPRESSED_READ  (97),
		.IN_PKT_BURSTWRAP_H            (109),
		.IN_PKT_BURSTWRAP_L            (107),
		.IN_PKT_BURST_SIZE_H           (112),
		.IN_PKT_BURST_SIZE_L           (110),
		.IN_PKT_RESPONSE_STATUS_H      (136),
		.IN_PKT_RESPONSE_STATUS_L      (135),
		.IN_PKT_TRANS_EXCLUSIVE        (102),
		.IN_PKT_BURST_TYPE_H           (114),
		.IN_PKT_BURST_TYPE_L           (113),
		.IN_ST_DATA_W                  (137),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (100),
		.OUT_PKT_RESPONSE_STATUS_L     (99),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (101),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (clk_50),                              //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_012_src_valid),             //      sink.valid
		.in_channel           (id_router_012_src_channel),           //          .channel
		.in_startofpacket     (id_router_012_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_012_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_012_src_ready),             //          .ready
		.in_data              (id_router_012_src_data),              //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_007_src_data),          //          .data
		.out_channel          (width_adapter_007_src_channel),       //          .channel
		.out_valid            (width_adapter_007_src_valid),         //          .valid
		.out_ready            (width_adapter_007_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	system_0_irq_mapper irq_mapper (
		.clk           (clk_50),                             //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (cpu_0_d_irq_irq)                     //    sender.irq
	);

endmodule
